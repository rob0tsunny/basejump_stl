module bsg_test_master
  #(
  )
  (
    input clk_i
    , input reset_i

    , input v_i
    , input write_not_read_i
    , input addr_i
  );


endmodule 
